`include "test_ldi.vh"
`include "test_in.vh"
`include "test_out.vh"
`include "test_sbi.vh"
`include "test_cbi.vh"
